module Half_adder(input a,b, output sum,carry);
{carry,sum} = a+b;
endmodule 
